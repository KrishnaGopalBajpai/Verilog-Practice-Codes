//AND gate using assign statement.


module andgt1 (f,a,b);
input a,b;
output f;
assign f=a&b;
enmodule
